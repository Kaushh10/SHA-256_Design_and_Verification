//A different approach to our Hashcore logic code
